package abc;
  class x;
      string q[$];
  endclass
endpackage

module sv_queue_example;
endmodule
