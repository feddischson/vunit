module string_example;


  function int example( string abc );

    if( abc[0] ) begin
      return 1;
    end else begin
      return 0;
    end

  endfunction


endmodule
