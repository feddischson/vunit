class top;
typedef enum 
{
X,
Y
} xy;
endclass
